module xor2 (A, B, Z);
    input A, B;
    output Z;
    
    xor(Z, A, B);
endmodule
